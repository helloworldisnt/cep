module sg13g2_Corner(); endmodule
